module test (

); 
endmodule