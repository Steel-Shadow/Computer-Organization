module mips (
    input clk,
    input reset
);
/************   declaration    ************/

/************   stage_F    ************/

/************   stage_D    ************/

/************   stage_E    ************/
/************   stage_M    ************/
/************   stage_W    ************/

endmodule
